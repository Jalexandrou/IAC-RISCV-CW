Test/ALU.sv