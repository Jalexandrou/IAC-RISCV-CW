module ALUDecoder #()(
    input [2:0] funct3,
    input [4:0] funct7,
    input logic op5,
    input [1:0] ALUOp
);

endmodule
