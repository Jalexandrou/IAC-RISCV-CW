module ALUDecoder #()(
    input  [2:0]    func3,
    input  [4:0]    func7,
    input  logic    op5,
    input  [1:0]    ALUOp,

    output [2:0]    ALUControl_o
);

endmodule
